/*
    mux主要功能是多路选择器。mux包含二选一、四选一多路选择器。
    信号名	方向	描述
    d0、d1、d2...	I	供选择数据（d0、d1）
    s	I	片选信号
    y	O	片选后的数据
*/
`timescale 1ns / 1ns
module MUX
        (
            input s;            //片选信号
            input y；           //片选后的数据
        );

        




endmodule