/*
    IMnoc是指令存储器，主要功能是根据读控制信号DMWr，读写对应addr地址的32位数据
    
    1	读指令存储器	输出地址所对应的指令，q imem[address]
*/
`timescale 1ns /  1ns
module IMnoc
			(
				input [9:0] address,   //访问地址
				output reg [31:0] dout     //读出的指令
			);

			//输出地址所对应的指令，q <- imem[address]
			reg [31:0] imem [0:31];
			initial begin
//				imem[0]=32'b00000000001000100001100000100011;//subu $1 $2 $3;
//				imem[1]=32'b00000000001000100001100000100001;//addu $1 $2 $3
//				imem[2]=32'b001101_00010_00001_0000000000000101;//ori $2 5 $1;
//				imem[3]=32'b101011_00001_10000_0000000000000001;//sw $16 1($1);
//				imem[4]=32'b001101_00000_10000_0000011111110011;//ori $16,$0, 11111110011;
//				imem[5]=32'b100011_00001_10000_0000000000000001;//lw $16 1($1);
////				imem[5]=32'b000100_00011_00000_1111111111111110;//beq $3 $0 -2;
////				imem[6]=32'b000100_00011_00011_1111111111111110;//beq $3 $3 -2;
////				imem[7]=32'b00001100_00000000_00001100_00000000;// jal 0x3000;

      //imem[0]=32'b000000_00001_00010_0001100000100011;
      //imem[1]=32'h0c000c01; // jal 0x3004
      
        imem[0]=32'b000000_00001_00010_0001100000100011;//subu $1 $2 $3
        imem[1]=32'b000000_00001_00010_0001100000100001;//addu $1 $2 $3
        imem[2]=32'b001101_00010_00001_0000000000000101;//ori $2 5 $1;
        imem[3]=32'b101011_00001_10000_0000000000000001;//sw $16 1($1);
        imem[4]=32'b001101_00000_10000_0000011111110011;//ori $16, $0, 11111110011;
        imem[5]=32'b100011_00001_10000_0000000000000001;//lw $16 1($1);
        
        
        imem[6]=32'h340b0000;// ori $11, $0, 0
        imem[7]=32'h340c0001;// ori $12, $0, 1
        imem[8]=32'h340d0001;// ori $13. $0, 1
        // the_loop: 0x00003009
        imem[9]=32'h016d5821;// addu $11, $11, $13
        imem[10]=32'h116cfffe;// beq $11, $12, the_loop
        imem[11]=32'h0c000c00;// jal 0x3000
		  
			end
			always@(*)begin
				dout = imem[address];
			end

endmodule